-- ========================================================
-- from VHDL producer:

-- Module ID: 2

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_0_1

-- Unique ID of L1 Trigger Menu:
-- 88611f82-f9d5-4db8-917c-95d140b6644a

-- Unique ID of firmware implementation:
-- c9eecec0-6ade-4733-b1f9-31711d57aa7c

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.13.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i113 : std_logic;
    signal single_ext_i139 : std_logic;
    signal single_ext_i86 : std_logic;
    signal single_ext_i91 : std_logic;
    signal single_htt_i112 : std_logic;
    signal single_eg_i118 : std_logic;
    signal single_jet_i119 : std_logic;
    signal single_jet_i125 : std_logic;
    signal single_jet_i126 : std_logic;
    signal single_mu_i129 : std_logic;
    signal single_mu_i133 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_beam_gas_b2_vme : std_logic;
    signal l1_bptx_or_ref4_vme : std_logic;
    signal l1_htt360er : std_logic;
    signal l1_last_collision_in_train : std_logic;
    signal l1_single_eg8er2p5 : std_logic;
    signal l1_single_jet120 : std_logic;
    signal l1_single_jet35_fwd3p0 : std_logic;
    signal l1_single_mu0_bmtf : std_logic;
    signal l1_single_mu22 : std_logic;
    signal l1_unpaired_bunch_bptx_plus : std_logic;

-- ========================================================