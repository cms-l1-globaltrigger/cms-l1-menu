-- ========================================================
-- from VHDL producer:

-- Module ID: 2

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2024_v1_0_5

-- Unique ID of L1 Trigger Menu:
-- 11642ab9-3cb5-4a4c-9431-46bf1ceb9bb7

-- Unique ID of firmware implementation:
-- 95dcc552-ab20-4c4f-8638-3b1c2079dbb4

-- Scale set:
-- scales_2023_02_16

-- VHDL producer
-- version: 2.20.1
-- hash value: 37aeed0f04da76b667e2567c8eee7fb6e0bbfdcc7e4a47a65d22d7168cf55357

-- tmEventSetup
-- version: 0.13.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i172 : std_logic;
    signal single_ext_i24 : std_logic;
    signal single_ext_i4 : std_logic;
    signal single_ext_i9 : std_logic;
    signal single_etmhf_i35 : std_logic;
    signal single_htt_i177 : std_logic;
    signal single_htt_i38 : std_logic;
    signal single_eg_i180 : std_logic;
    signal single_eg_i185 : std_logic;
    signal single_eg_i252 : std_logic;
    signal single_eg_i256 : std_logic;
    signal single_jet_i187 : std_logic;
    signal single_jet_i51 : std_logic;
    signal single_jet_i54 : std_logic;
    signal single_jet_i55 : std_logic;
    signal single_jet_i56 : std_logic;
    signal single_mu_i59 : std_logic;
    signal single_mu_i60 : std_logic;
    signal single_mu_i61 : std_logic;
    signal triple_eg_i199 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_beam_gas_b1_vme : std_logic;
    signal l1_bptx_or_ref3_vme : std_logic;
    signal l1_unpaired_bunch_bptx_plus : std_logic;
    signal l1_etmhf100 : std_logic;
    signal l1_htt200er : std_logic;
    signal l1_htt400er : std_logic;
    signal l1_hcal_laser_mon_trig : std_logic;
    signal l1_single_eg34er2p5 : std_logic;
    signal l1_single_eg45er2p5 : std_logic;
    signal l1_triple_eg_18_17_8_er2p5 : std_logic;
    signal l1_single_jet8er_he : std_logic;
    signal l1_single_jet35er2p5 : std_logic;
    signal l1_single_jet120 : std_logic;
    signal l1_single_jet120_fwd3p0 : std_logic;
    signal l1_single_mu0_dq : std_logic;
    signal l1_single_mu0_bmtf : std_logic;
    signal l1_single_mu0_emtf : std_logic;
    signal l1_single_mu22_emtf : std_logic;
    signal l1_single_iso_eg26er2p1 : std_logic;
    signal l1_single_iso_eg30er2p1 : std_logic;

-- ========================================================