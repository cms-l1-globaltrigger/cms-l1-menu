-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2024_v1_0_5

-- Unique ID of L1 Trigger Menu:
-- 11642ab9-3cb5-4a4c-9431-46bf1ceb9bb7

-- Unique ID of firmware implementation:
-- 95dcc552-ab20-4c4f-8638-3b1c2079dbb4

-- Scale set:
-- scales_2023_02_16

-- VHDL producer
-- version: 2.20.1
-- hash value: 37aeed0f04da76b667e2567c8eee7fb6e0bbfdcc7e4a47a65d22d7168cf55357

-- tmEventSetup
-- version: 0.13.0

-- Signal definition of pt, eta and phi for correlation conditions.
    signal tau_bx_0_pt_vector: diff_inputs_array(0 to NR_TAU_OBJECTS-1) := (others => (others => '0'));
    signal tau_bx_0_eta_integer: integer_array(0 to NR_TAU_OBJECTS-1) := (others => 0);
    signal tau_bx_0_phi_integer: integer_array(0 to NR_TAU_OBJECTS-1) := (others => 0);
    signal tau_bx_0_cos_phi: integer_array(0 to NR_TAU_OBJECTS-1) := (others => 0);
    signal tau_bx_0_sin_phi: integer_array(0 to NR_TAU_OBJECTS-1) := (others => 0);
    signal tau_bx_0_conv_cos_phi: integer_array(0 to NR_TAU_OBJECTS-1) := (others => 0);
    signal tau_bx_0_conv_sin_phi: integer_array(0 to NR_TAU_OBJECTS-1) := (others => 0);
    signal tau_bx_0_eta_conv_2_muon_eta_integer: integer_array(0 to NR_TAU_OBJECTS-1) := (others => 0);
    signal tau_bx_0_phi_conv_2_muon_phi_integer: integer_array(0 to NR_TAU_OBJECTS-1) := (others => 0);
    signal jet_bx_0_pt_vector: diff_inputs_array(0 to NR_JET_OBJECTS-1) := (others => (others => '0'));
    signal jet_bx_0_eta_integer: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_phi_integer: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_cos_phi: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_sin_phi: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_conv_cos_phi: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_conv_sin_phi: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_eta_conv_2_muon_eta_integer: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_phi_conv_2_muon_phi_integer: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal mu_bx_0_pt_vector: diff_inputs_array(0 to NR_MU_OBJECTS-1) := (others => (others => '0'));
    signal mu_bx_0_upt_vector: diff_inputs_array(0 to NR_MU_OBJECTS-1) := (others => (others => '0'));
    signal mu_bx_0_eta_integer: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_phi_integer: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_eta_integer_half_res: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_phi_integer_half_res: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_cos_phi: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_sin_phi: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);

-- Signal definition for cuts of correlation conditions.
    signal tau_tau_bx_0_bx_0_deta_integer: dim2_max_eta_range_array(0 to NR_TAU_OBJECTS-1, 0 to NR_TAU_OBJECTS-1) := (others => (others => 0));
    signal tau_tau_bx_0_bx_0_deta: deta_dphi_vector_array(0 to NR_TAU_OBJECTS-1, 0 to NR_TAU_OBJECTS-1) := (others => (others => (others => '0')));
    signal tau_tau_bx_0_bx_0_dphi_integer: dim2_max_phi_range_array(0 to NR_TAU_OBJECTS-1, 0 to NR_TAU_OBJECTS-1) := (others => (others => 0));
    signal tau_tau_bx_0_bx_0_dphi: deta_dphi_vector_array(0 to NR_TAU_OBJECTS-1, 0 to NR_TAU_OBJECTS-1) := (others => (others => (others => '0')));
    signal jet_jet_bx_0_bx_0_deta_integer: dim2_max_eta_range_array(0 to NR_JET_OBJECTS-1, 0 to NR_JET_OBJECTS-1) := (others => (others => 0));
    signal jet_jet_bx_0_bx_0_deta: deta_dphi_vector_array(0 to NR_JET_OBJECTS-1, 0 to NR_JET_OBJECTS-1) := (others => (others => (others => '0')));
    signal jet_jet_bx_0_bx_0_dphi_integer: dim2_max_phi_range_array(0 to NR_JET_OBJECTS-1, 0 to NR_JET_OBJECTS-1) := (others => (others => 0));
    signal jet_jet_bx_0_bx_0_dphi: deta_dphi_vector_array(0 to NR_JET_OBJECTS-1, 0 to NR_JET_OBJECTS-1) := (others => (others => (others => '0')));
    signal mu_mu_bx_0_bx_0_deta_integer: dim2_max_eta_range_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => 0));
    signal mu_mu_bx_0_bx_0_deta: deta_dphi_vector_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => (others => '0')));
    signal mu_mu_bx_0_bx_0_dphi_integer: dim2_max_phi_range_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => 0));
    signal mu_mu_bx_0_bx_0_dphi: deta_dphi_vector_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => (others => '0')));
    signal mu_mu_bx_0_bx_0_deta_integer_half_res: dim2_max_eta_range_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => 0));
    signal mu_mu_bx_0_bx_0_dphi_integer_half_res: dim2_max_phi_range_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => 0));
    signal mu_mu_bx_0_bx_0_dr : dr_dim2_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => (others => '0')));
    signal mu_mu_bx_0_bx_0_mass_inv_pt : mass_dim2_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => (others => '0')));

-- Signal definition for muon charge correlations.
    signal ls_charcorr_double_bx_0_bx_0, os_charcorr_double_bx_0_bx_0 : std_logic_2dim_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1);
    signal ls_charcorr_triple_bx_0_bx_0, os_charcorr_triple_bx_0_bx_0 : std_logic_3dim_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1);
    signal ls_charcorr_quad_bx_0_bx_0, os_charcorr_quad_bx_0_bx_0 : std_logic_4dim_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1);

-- Signal definition for conditions names
    signal single_cent0_i28 : std_logic;
    signal single_cent1_i29 : std_logic;
    signal single_cent2_i30 : std_logic;
    signal single_cent3_i31 : std_logic;
    signal single_cent4_i32 : std_logic;
    signal single_cent5_i140 : std_logic;
    signal single_cent6_i139 : std_logic;
    signal single_cent7_i201 : std_logic;
    signal single_ext_i0 : std_logic;
    signal single_ext_i14 : std_logic;
    signal single_ext_i15 : std_logic;
    signal single_ext_i16 : std_logic;
    signal single_ext_i17 : std_logic;
    signal single_ext_i18 : std_logic;
    signal single_ext_i19 : std_logic;
    signal single_ext_i20 : std_logic;
    signal single_ext_i21 : std_logic;
    signal single_ext_i22 : std_logic;
    signal single_ext_i27 : std_logic;
    signal single_mbt0_hfm_i34 : std_logic;
    signal single_mbt1_hfm_i131 : std_logic;
    signal single_mbt0_hfp_i33 : std_logic;
    signal single_mbt1_hfp_i130 : std_logic;
    signal muon_shower0_i142 : std_logic;
    signal muon_shower1_i141 : std_logic;
    signal single_towercount_i240 : std_logic;
    signal zdc_minus_i135 : std_logic;
    signal zdc_minus_i144 : std_logic;
    signal zdc_minus_i146 : std_logic;
    signal zdc_minus_i148 : std_logic;
    signal zdc_minus_i151 : std_logic;
    signal zdc_minus_i153 : std_logic;
    signal zdc_minus_i155 : std_logic;
    signal zdc_minus_i157 : std_logic;
    signal zdc_minus_i159 : std_logic;
    signal zdc_minus_i161 : std_logic;
    signal zdc_minus_i163 : std_logic;
    signal zdc_minus_i206 : std_logic;
    signal zdc_minus_i237 : std_logic;
    signal zdc_minus_i238 : std_logic;
    signal zdc_minus_i248 : std_logic;
    signal zdc_minus_i250 : std_logic;
    signal zdc_plus_i134 : std_logic;
    signal zdc_plus_i143 : std_logic;
    signal zdc_plus_i145 : std_logic;
    signal zdc_plus_i147 : std_logic;
    signal zdc_plus_i150 : std_logic;
    signal zdc_plus_i152 : std_logic;
    signal zdc_plus_i154 : std_logic;
    signal zdc_plus_i156 : std_logic;
    signal zdc_plus_i158 : std_logic;
    signal zdc_plus_i160 : std_logic;
    signal zdc_plus_i162 : std_logic;
    signal zdc_plus_i207 : std_logic;
    signal zdc_plus_i236 : std_logic;
    signal zdc_plus_i239 : std_logic;
    signal zdc_plus_i247 : std_logic;
    signal zdc_plus_i249 : std_logic;
    signal calo_calo_correlation_i230 : std_logic;
    signal calo_calo_correlation_i231 : std_logic;
    signal calo_calo_correlation_i232 : std_logic;
    signal calo_calo_correlation_i233 : std_logic;
    signal calo_calo_correlation_i234 : std_logic;
    signal calo_calo_correlation_i235 : std_logic;
    signal calo_calo_correlation_i244 : std_logic;
    signal calo_calo_correlation_i245 : std_logic;
    signal calo_calo_correlation_i246 : std_logic;
    signal invariant_mass_i117 : std_logic;
    signal invariant_mass_i118 : std_logic;
    signal invariant_mass_i119 : std_logic;
    signal muon_muon_correlation_i114 : std_logic;
    signal muon_muon_correlation_i115 : std_logic;
    signal muon_muon_correlation_i116 : std_logic;
    signal double_eg_i100 : std_logic;
    signal double_eg_i101 : std_logic;
    signal double_eg_i136 : std_logic;
    signal double_eg_i137 : std_logic;
    signal double_eg_i98 : std_logic;
    signal double_eg_i99 : std_logic;
    signal double_mu_i109 : std_logic;
    signal double_mu_i110 : std_logic;
    signal double_mu_i111 : std_logic;
    signal double_mu_i112 : std_logic;
    signal double_mu_i113 : std_logic;
    signal double_mu_i133 : std_logic;
    signal double_mu_i67 : std_logic;
    signal single_eg_i102 : std_logic;
    signal single_eg_i103 : std_logic;
    signal single_eg_i126 : std_logic;
    signal single_eg_i127 : std_logic;
    signal single_eg_i128 : std_logic;
    signal single_eg_i138 : std_logic;
    signal single_eg_i202 : std_logic;
    signal single_eg_i41 : std_logic;
    signal single_eg_i42 : std_logic;
    signal single_eg_i96 : std_logic;
    signal single_eg_i97 : std_logic;
    signal single_jet_i120 : std_logic;
    signal single_jet_i121 : std_logic;
    signal single_jet_i122 : std_logic;
    signal single_jet_i123 : std_logic;
    signal single_jet_i124 : std_logic;
    signal single_jet_i125 : std_logic;
    signal single_jet_i149 : std_logic;
    signal single_jet_i205 : std_logic;
    signal single_jet_i208 : std_logic;
    signal single_jet_i209 : std_logic;
    signal single_jet_i210 : std_logic;
    signal single_jet_i211 : std_logic;
    signal single_jet_i212 : std_logic;
    signal single_jet_i213 : std_logic;
    signal single_jet_i214 : std_logic;
    signal single_jet_i215 : std_logic;
    signal single_jet_i216 : std_logic;
    signal single_jet_i217 : std_logic;
    signal single_jet_i218 : std_logic;
    signal single_jet_i219 : std_logic;
    signal single_jet_i241 : std_logic;
    signal single_jet_i242 : std_logic;
    signal single_jet_i243 : std_logic;
    signal single_jet_i52 : std_logic;
    signal single_jet_i69 : std_logic;
    signal single_jet_i70 : std_logic;
    signal single_jet_i71 : std_logic;
    signal single_jet_i72 : std_logic;
    signal single_jet_i73 : std_logic;
    signal single_jet_i74 : std_logic;
    signal single_jet_i75 : std_logic;
    signal single_jet_i76 : std_logic;
    signal single_jet_i77 : std_logic;
    signal single_jet_i78 : std_logic;
    signal single_jet_i79 : std_logic;
    signal single_jet_i80 : std_logic;
    signal single_jet_i81 : std_logic;
    signal single_jet_i82 : std_logic;
    signal single_jet_i83 : std_logic;
    signal single_jet_i84 : std_logic;
    signal single_jet_i85 : std_logic;
    signal single_jet_i86 : std_logic;
    signal single_jet_i87 : std_logic;
    signal single_jet_i88 : std_logic;
    signal single_jet_i89 : std_logic;
    signal single_jet_i90 : std_logic;
    signal single_jet_i91 : std_logic;
    signal single_jet_i92 : std_logic;
    signal single_jet_i93 : std_logic;
    signal single_jet_i94 : std_logic;
    signal single_jet_i95 : std_logic;
    signal single_mu_i104 : std_logic;
    signal single_mu_i105 : std_logic;
    signal single_mu_i106 : std_logic;
    signal single_mu_i107 : std_logic;
    signal single_mu_i108 : std_logic;
    signal single_mu_i129 : std_logic;
    signal single_mu_i132 : std_logic;
    signal single_mu_i193 : std_logic;
    signal single_mu_i194 : std_logic;
    signal single_mu_i229 : std_logic;
    signal single_mu_i66 : std_logic;
    signal single_tau_i220 : std_logic;
    signal single_tau_i221 : std_logic;
    signal single_tau_i222 : std_logic;
    signal single_tau_i223 : std_logic;
    signal single_tau_i224 : std_logic;
    signal single_tau_i225 : std_logic;
    signal single_tau_i226 : std_logic;
    signal single_tau_i227 : std_logic;
    signal single_tau_i228 : std_logic;

-- Signal definition for algorithms names
    signal l1_always_true : std_logic;
    signal l1_zero_bias : std_logic;
    signal l1_zero_bias_copy : std_logic;
    signal l1_bptx_or : std_logic;
    signal l1_not_bptx_or : std_logic;
    signal l1_first_bunch_after_train : std_logic;
    signal l1_first_bunch_before_train : std_logic;
    signal l1_first_bunch_in_train : std_logic;
    signal l1_isolated_bunch : std_logic;
    signal l1_last_bunch_in_train : std_logic;
    signal l1_second_bunch_in_train : std_logic;
    signal l1_second_last_bunch_in_train : std_logic;
    signal l1_first_collision_in_orbit : std_logic;
    signal l1_first_collision_in_orbit_centrality30_100_bptx_and : std_logic;
    signal l1_first_collision_in_orbit_centrality50_100_bptx_and : std_logic;
    signal l1_single_eg3 : std_logic;
    signal l1_single_eg5 : std_logic;
    signal l1_minimum_bias_hf1_and_bptx_and_copy : std_logic;
    signal l1_zdc1n_or_minimum_bias_hf1_and_bptx_and_copy : std_logic;
    signal l1_zdc2n_or_minimum_bias_hf1_and_bptx_and_copy : std_logic;
    signal l1_single_jet60 : std_logic;
    signal l1_single_mu_open : std_logic;
    signal l1_single_mu_open_not_bptx_or : std_logic;
    signal l1_single_mu_open_er1p4_not_bptx_or_3_bx : std_logic;
    signal l1_single_mu_open_er1p1_not_bptx_or_3_bx : std_logic;
    signal l1_single_mu_cosmics : std_logic;
    signal l1_single_mu_cosmics_emtf : std_logic;
    signal l1_single_mu3 : std_logic;
    signal l1_single_mu5 : std_logic;
    signal l1_single_mu7 : std_logic;
    signal l1_double_mu0 : std_logic;
    signal l1_double_mu0_sq : std_logic;
    signal l1_single_mu_open_centrality_30_100_bptx_and : std_logic;
    signal l1_single_mu0_centrality_40_100_bptx_and : std_logic;
    signal l1_single_mu0_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet28_bptx_and : std_logic;
    signal l1_single_jet28_d_meson_bptx_and : std_logic;
    signal l1_single_jet32_bptx_and : std_logic;
    signal l1_single_jet36_bptx_and : std_logic;
    signal l1_single_jet40_bptx_and : std_logic;
    signal l1_single_jet44_bptx_and : std_logic;
    signal l1_single_jet44_d_meson_bptx_and : std_logic;
    signal l1_single_jet48_bptx_and : std_logic;
    signal l1_single_jet56_bptx_and : std_logic;
    signal l1_single_jet60_bptx_and : std_logic;
    signal l1_single_jet60_d_meson_bptx_and : std_logic;
    signal l1_single_jet64_bptx_and : std_logic;
    signal l1_single_jet72_bptx_and : std_logic;
    signal l1_single_jet80_bptx_and : std_logic;
    signal l1_single_jet8_fwd_bptx_and : std_logic;
    signal l1_single_jet16_fwd_bptx_and : std_logic;
    signal l1_single_jet28_fwd_bptx_and : std_logic;
    signal l1_single_jet36_fwd_bptx_and : std_logic;
    signal l1_single_jet44_fwd_bptx_and : std_logic;
    signal l1_single_jet56_fwd_bptx_and : std_logic;
    signal l1_single_jet64_fwd_bptx_and : std_logic;
    signal l1_single_jet8_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet16_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet24_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet28_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet32_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet36_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet40_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet44_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet48_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet56_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet60_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet64_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet8_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet16_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet24_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet28_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet32_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet36_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet40_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet44_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet48_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet56_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet60_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet64_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet8_bptx_and : std_logic;
    signal l1_single_jet16_bptx_and : std_logic;
    signal l1_single_jet24_bptx_and : std_logic;
    signal l1_double_mu0_sq_bptx_and : std_logic;
    signal l1_single_eg3_bptx_and : std_logic;
    signal l1_single_eg4_bptx_and : std_logic;
    signal l1_single_eg5_bptx_and : std_logic;
    signal l1_single_eg7_bptx_and : std_logic;
    signal l1_single_eg12_bptx_and : std_logic;
    signal l1_single_eg15_bptx_and : std_logic;
    signal l1_single_eg21_bptx_and : std_logic;
    signal l1_single_eg30_bptx_and : std_logic;
    signal l1_double_eg2_bptx_and : std_logic;
    signal l1_double_eg5_bptx_and : std_logic;
    signal l1_double_eg8_bptx_and : std_logic;
    signal l1_double_eg10_bptx_and : std_logic;
    signal l1_single_eg3_centrality_30_100_bptx_and : std_logic;
    signal l1_single_eg7_centrality_30_100_bptx_and : std_logic;
    signal l1_single_eg15_centrality_30_100_bptx_and : std_logic;
    signal l1_single_eg21_centrality_30_100_bptx_and : std_logic;
    signal l1_single_mu_open_bptx_and : std_logic;
    signal l1_single_mu3_open_bptx_and : std_logic;
    signal l1_single_mu0_bptx_and : std_logic;
    signal l1_single_mu3_bptx_and : std_logic;
    signal l1_single_mu5_bptx_and : std_logic;
    signal l1_single_mu7_bptx_and : std_logic;
    signal l1_double_mu_open_bptx_and : std_logic;
    signal l1_double_mu_open_os_bptx_and : std_logic;
    signal l1_double_mu_open_ss_bptx_and : std_logic;
    signal l1_double_mu_open_max_dr3p5_bptx_and : std_logic;
    signal l1_double_mu_open_max_dr3p5_m0to7_bptx_and : std_logic;
    signal l1_double_mu_sq_bptx_and : std_logic;
    signal l1_double_mu_sq_max_dr3p5_bptx_and : std_logic;
    signal l1_double_mu_sq_max_dr3p5_m0to7_bptx_and : std_logic;
    signal l1_double_mu0_bptx_and : std_logic;
    signal l1_double_mu0_max_dr3p5_bptx_and : std_logic;
    signal l1_double_mu0_max_dr3p5_m0to7_bptx_and : std_logic;
    signal l1_double_mu10_bptx_and : std_logic;
    signal l1_double_mu_open_centrality_30_100_bptx_and : std_logic;
    signal l1_double_mu_open_centrality_40_100_bptx_and : std_logic;
    signal l1_double_mu_open_centrality_50_100_bptx_and : std_logic;
    signal l1_single_mu_open_single_jet28_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu_open_single_jet44_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu_open_single_jet56_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu_open_single_jet64_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu3_single_jet28_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu3_single_jet32_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu3_single_jet40_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu_open_single_eg15_bptx_and : std_logic;
    signal l1_single_mu3_single_eg12_bptx_and : std_logic;
    signal l1_single_mu3_single_eg20_bptx_and : std_logic;
    signal l1_single_mu3_single_eg30_bptx_and : std_logic;
    signal l1_single_mu5_single_eg10_bptx_and : std_logic;
    signal l1_single_mu5_single_eg12_bptx_and : std_logic;
    signal l1_single_mu5_single_eg15_bptx_and : std_logic;
    signal l1_single_mu5_single_eg20_bptx_and : std_logic;
    signal l1_single_mu7_single_eg7_bptx_and : std_logic;
    signal l1_single_mu7_single_eg10_bptx_and : std_logic;
    signal l1_single_mu7_single_eg12_bptx_and : std_logic;
    signal l1_single_mu7_single_eg15_bptx_and : std_logic;
    signal l1_single_mu12_single_eg7_bptx_and : std_logic;
    signal l1_single_mu_cosmic_bptx_and : std_logic;
    signal l1_single_mu_cosmic_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_mu_cosmic_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_mu_cosmic_bptx_and : std_logic;
    signal l1_double_mu_cosmic_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_mu_open_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_mu_open_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_mu_open_or_single_mu_cosmic_emtf_bptx_and : std_logic;
    signal l1_single_mu_open_or_single_mu_cosmic_emtf_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_mu_open_or_single_mu_cosmic_emtf_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_mu_open_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_mu0_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_eg3_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_eg4_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_eg2_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_eg3_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_eg4_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_eg5_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_eg1_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_eg2_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_eg3_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_eg5_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_mu_shower_tight : std_logic;
    signal l1_single_mu_shower_nominal : std_logic;
    signal l1_single_mu_shower_tight_bptx_and : std_logic;
    signal l1_single_mu_shower_nominal_bptx_and : std_logic;
    signal l1_centrality_saturation_bptx_and : std_logic;
    signal l1_centrality_0_0p5_bptx_and : std_logic;
    signal l1_centrality_0_1_bptx_and : std_logic;
    signal l1_centrality_30_40_bptx_and : std_logic;
    signal l1_centrality_40_50_bptx_and : std_logic;
    signal l1_centrality_30_50_bptx_and : std_logic;
    signal l1_centrality_50_65_bptx_and : std_logic;
    signal l1_centrality_65_80_bptx_and : std_logic;
    signal l1_centrality_80_100_bptx_and : std_logic;
    signal l1_centrality_30_100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_centrality_50_100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_zdc1n_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp1_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp2_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp3_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc2n_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc2n_bkp1_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc2n_bkp2_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc2n_bkp3_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc3n_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc3n_bkp1_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc3n_bkp2_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc3n_bkp3_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_and_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp1_and_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp2_and_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp3_and_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_zdc1n_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp1_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp2_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp3_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc2n_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc2n_bkp1_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc2n_bkp2_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc2n_bkp3_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc3n_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc3n_bkp1_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc3n_bkp2_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc3n_bkp3_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_and_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp1_and_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp2_and_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp3_and_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_eg2_zdc1n_or_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_or_bptx_and : std_logic;
    signal l1_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_zdc1n_xor_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp1_xor_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp2_xor_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp3_xor_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_asym_xor_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp1_asym_xor_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp2_asym_xor_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_xor_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp1_xor_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp2_xor_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_asym_xor_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp1_asym_xor_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp2_asym_xor_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_jet8_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_jet8_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_jet12_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_jet12_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_jet16_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_jet16_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_jet20_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_jet20_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_jet24_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_jet24_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_jet28_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_jet28_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_jet8_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_jet12_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_jet16_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_jet20_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_jet24_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_jet28_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdcp14 : std_logic;
    signal l1_zdcp14_bptx_and : std_logic;
    signal l1_zdcm14 : std_logic;
    signal l1_zdcm14_bptx_and : std_logic;
    signal l1_zdc14_and : std_logic;
    signal l1_zdc14_and_bptx_and : std_logic;
    signal l1_zdc14_or : std_logic;
    signal l1_zdc14_or_bptx_and : std_logic;
    signal l1_zdcp16 : std_logic;
    signal l1_zdcp16_bptx_and : std_logic;
    signal l1_zdcm16 : std_logic;
    signal l1_zdcm16_bptx_and : std_logic;
    signal l1_zdc16_and : std_logic;
    signal l1_zdc16_and_bptx_and : std_logic;
    signal l1_zdc16_or : std_logic;
    signal l1_zdc16_or_bptx_and : std_logic;
    signal l1_zdcp18 : std_logic;
    signal l1_zdcp18_bptx_and : std_logic;
    signal l1_zdcm18 : std_logic;
    signal l1_zdcm18_bptx_and : std_logic;
    signal l1_zdc18_and : std_logic;
    signal l1_zdc18_and_bptx_and : std_logic;
    signal l1_zdc18_or : std_logic;
    signal l1_zdc18_or_bptx_and : std_logic;
    signal l1_zdcp22 : std_logic;
    signal l1_zdcp22_bptx_and : std_logic;
    signal l1_zdcm22 : std_logic;
    signal l1_zdcm22_bptx_and : std_logic;
    signal l1_zdc22_and : std_logic;
    signal l1_zdc22_and_bptx_and : std_logic;
    signal l1_zdc22_or : std_logic;
    signal l1_zdc22_or_bptx_and : std_logic;
    signal l1_zdcp28 : std_logic;
    signal l1_zdcp28_bptx_and : std_logic;
    signal l1_zdcm28 : std_logic;
    signal l1_zdcm28_bptx_and : std_logic;
    signal l1_zdc28_and : std_logic;
    signal l1_zdc28_and_bptx_and : std_logic;
    signal l1_zdc28_or : std_logic;
    signal l1_zdc28_or_bptx_and : std_logic;
    signal l1_zdc1n_and_and_not_mbhf2_bptx_and : std_logic;
    signal l1_zdc1n_and_and_not_mbhf2_or_bptx_and : std_logic;
    signal l1_single_jet8_zdc1n_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet8_zdc1n_asym_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet12_zdc1n_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet12_zdc1n_asym_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet16_zdc1n_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet16_zdc1n_asym_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet20_zdc1n_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet20_zdc1n_asym_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet24_zdc1n_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet24_zdc1n_asym_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet28_zdc1n_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_jet28_zdc1n_asym_xor_not_pre_bptx_bptx_and : std_logic;
    signal l1_single_uncorr_jet2_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet4_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet6_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet8_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet12_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet16_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet20_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet24_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet28_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp3_asym_xor_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp3_xor_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc1n_bkp3_asym_xor_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet2_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet4_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet6_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet8_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet12_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet16_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet20_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet24_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet28_zdc1n_bkp1_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet2_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet4_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet6_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet8_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet12_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet16_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet20_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet24_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet28_zdc1n_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet2_zdc1n_bkp1_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet4_zdc1n_bkp1_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet6_zdc1n_bkp1_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet8_zdc1n_bkp1_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet12_zdc1n_bkp1_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet16_zdc1n_bkp1_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet20_zdc1n_bkp1_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet24_zdc1n_bkp1_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet28_zdc1n_bkp1_xor_bptx_and : std_logic;
    signal l1_double_jet8_delta_phi2p0_not_zdc_or_bptx_and : std_logic;
    signal l1_double_jet12_delta_phi2p0_not_zdc_or_bptx_and : std_logic;
    signal l1_double_jet16_delta_phi2p0_not_zdc_or_bptx_and : std_logic;
    signal l1_double_uncorr_jet8_delta_phi2p0_not_zdc_or_bptx_and : std_logic;
    signal l1_double_uncorr_jet12_delta_phi2p0_not_zdc_or_bptx_and : std_logic;
    signal l1_double_uncorr_jet16_delta_phi2p0_not_zdc_or_bptx_and : std_logic;
    signal l1_double_jet8_delta_phi2p0_not_zdc1n_and_bptx_and : std_logic;
    signal l1_double_jet12_delta_phi2p0_not_zdc1n_and_bptx_and : std_logic;
    signal l1_double_jet16_delta_phi2p0_not_zdc1n_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet2_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet4_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet6_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet8_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet12_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet16_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet20_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet24_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet28_zdc1n_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet2_zdc1n_bkp1_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet4_zdc1n_bkp1_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet6_zdc1n_bkp1_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet8_zdc1n_bkp1_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet12_zdc1n_bkp1_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet16_zdc1n_bkp1_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet20_zdc1n_bkp1_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet24_zdc1n_bkp1_asym_xor_bptx_and : std_logic;
    signal l1_single_uncorr_jet28_zdc1n_bkp1_asym_xor_bptx_and : std_logic;
    signal l1_double_uncorr_jet2_delta_phi2p0_not_minimum_bias_hf2_bptx_and : std_logic;
    signal l1_double_uncorr_jet4_delta_phi2p0_not_minimum_bias_hf2_bptx_and : std_logic;
    signal l1_double_uncorr_jet6_delta_phi2p0_not_minimum_bias_hf2_bptx_and : std_logic;
    signal l1_double_uncorr_jet8_delta_phi2p0_not_minimum_bias_hf2_bptx_and : std_logic;
    signal l1_double_uncorr_jet12_delta_phi2p0_not_minimum_bias_hf2_bptx_and : std_logic;
    signal l1_double_uncorr_jet16_delta_phi2p0_not_minimum_bias_hf2_bptx_and : std_logic;
    signal l1_double_jet8_delta_phi2p0_not_minimum_bias_hf2_bptx_and : std_logic;
    signal l1_double_jet12_delta_phi2p0_not_minimum_bias_hf2_bptx_and : std_logic;
    signal l1_double_jet16_delta_phi2p0_not_minimum_bias_hf2_bptx_and : std_logic;
    signal l1_double_uncorr_jet2_delta_phi2p0_not_zdc1n_and_bptx_and : std_logic;
    signal l1_double_uncorr_jet4_delta_phi2p0_not_zdc1n_and_bptx_and : std_logic;
    signal l1_double_uncorr_jet6_delta_phi2p0_not_zdc1n_and_bptx_and : std_logic;
    signal l1_double_uncorr_jet8_delta_phi2p0_not_zdc1n_and_bptx_and : std_logic;
    signal l1_double_uncorr_jet12_delta_phi2p0_not_zdc1n_and_bptx_and : std_logic;
    signal l1_double_uncorr_jet16_delta_phi2p0_not_zdc1n_and_bptx_and : std_logic;
    signal l1_single_uncorr_jet2_not_zdc_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet4_not_zdc_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet6_not_zdc_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet8_not_zdc_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet12_not_zdc_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet16_not_zdc_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet20_not_zdc_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet24_not_zdc_or_bptx_and : std_logic;
    signal l1_single_uncorr_jet28_not_zdc_or_bptx_and : std_logic;
    signal l1_single_jet8_not_zdc_or_bptx_and : std_logic;
    signal l1_single_jet12_not_zdc_or_bptx_and : std_logic;
    signal l1_single_jet16_not_zdc_or_bptx_and : std_logic;
    signal l1_single_jet20_not_zdc_or_bptx_and : std_logic;
    signal l1_single_jet24_not_zdc_or_bptx_and : std_logic;
    signal l1_single_jet28_not_zdc_or_bptx_and : std_logic;
    signal l1_first_bunch_in_train_50ns : std_logic;
    signal l1_last_bunch_in_train_50ns : std_logic;
    signal l1_zdc1n_or_rap_gap_bptx_and : std_logic;
    signal l1_single_jet2_zdc1n_xor_rap_gap_bptx_and : std_logic;
    signal l1_single_jet4_zdc1n_xor_rap_gap_bptx_and : std_logic;
    signal l1_single_jet6_zdc1n_xor_rap_gap_bptx_and : std_logic;
    signal l1_single_jet8_zdc1n_xor_rap_gap_bptx_and : std_logic;
    signal l1_single_jet12_zdc1n_xor_rap_gap_bptx_and : std_logic;
    signal l1_single_jet16_zdc1n_xor_rap_gap_bptx_and : std_logic;
    signal l1_single_jet20_zdc1n_xor_rap_gap_bptx_and : std_logic;
    signal l1_single_jet24_zdc1n_xor_rap_gap_bptx_and : std_logic;
    signal l1_single_jet28_zdc1n_xor_rap_gap_bptx_and : std_logic;

-- ========================================================