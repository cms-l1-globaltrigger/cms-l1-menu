-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_1_0

-- Unique ID of L1 Trigger Menu:
-- 11f4244d-31e8-434f-b121-3188fa41b985

-- Unique ID of firmware implementation:
-- c8183b8a-5519-47a4-ad38-1ceb98bede21

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.13.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i82 : std_logic;
    signal single_ext_i87 : std_logic;
    signal single_ext_i92 : std_logic;
    signal muon_shower1_i59 : std_logic;
    signal single_ett_i98 : std_logic;
    signal single_jet_i122 : std_logic;
    signal single_jet_i124 : std_logic;
    signal single_mu_i131 : std_logic;
    signal single_mu_i134 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_and_ref1_vme : std_logic;
    signal l1_bptx_beam_gas_ref1_vme : std_logic;
    signal l1_bptx_ref_and_vme : std_logic;
    signal l1_mu_shower_one_tight : std_logic;
    signal l1_ett2000 : std_logic;
    signal l1_single_jet120er2p5 : std_logic;
    signal l1_single_jet35 : std_logic;
    signal l1_single_mu0_emtf : std_logic;
    signal l1_single_mu22_bmtf : std_logic;
    signal l1_single_mu22_emtf : std_logic;

-- ========================================================