-- ========================================================
-- from VHDL producer:

-- Module ID: 5

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_0_1

-- Unique ID of L1 Trigger Menu:
-- 88611f82-f9d5-4db8-917c-95d140b6644a

-- Unique ID of firmware implementation:
-- c9eecec0-6ade-4733-b1f9-31711d57aa7c

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.13.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i83 : std_logic;
    signal single_ext_i88 : std_logic;
    signal single_ext_i93 : std_logic;
    signal single_ext_i94 : std_logic;
    signal single_htt_i109 : std_logic;
    signal single_eg_i115 : std_logic;
    signal single_eg_i117 : std_logic;
    signal single_jet_i128 : std_logic;
    signal single_mu_i135 : std_logic;
    signal single_mu_i137 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_and_ref3_vme : std_logic;
    signal l1_bptx_beam_gas_ref2_vme : std_logic;
    signal l1_bptx_minus : std_logic;
    signal l1_bptx_minus_not_bptx_plus : std_logic;
    signal l1_bptx_plus : std_logic;
    signal l1_bptx_plus_not_bptx_minus : std_logic;
    signal l1_bptx_xor : std_logic;
    signal l1_htt120er : std_logic;
    signal l1_single_eg15er2p5 : std_logic;
    signal l1_single_eg50 : std_logic;
    signal l1_single_jet90 : std_logic;
    signal l1_single_mu22_omtf : std_logic;
    signal l1_single_mu_cosmics_omtf : std_logic;

-- ========================================================