-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2023_v0_0_3

-- Unique ID of L1 Trigger Menu:
-- 3caede45-ba4f-4464-8773-8dd386d7d3c4

-- Unique ID of firmware implementation:
-- 64f242dd-0bd3-48bc-aaed-b19fb8b7a2f3

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.14.2

-- tmEventSetup version
-- v0.11.2

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i1 : std_logic;
    signal single_ext_i11 : std_logic;
    signal single_ext_i24 : std_logic;
    signal single_ext_i6 : std_logic;
    signal single_ett_i36 : std_logic;
    signal single_jet_i48 : std_logic;
    signal single_jet_i57 : std_logic;
    signal single_mu_i61 : std_logic;
    signal single_mu_i64 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_and_ref1_vme : std_logic;
    signal l1_bptx_beam_gas_ref1_vme : std_logic;
    signal l1_bptx_ref_and_vme : std_logic;
    signal l1_unpaired_bunch_bptx_plus : std_logic;
    signal l1_ett2000 : std_logic;
    signal l1_single_jet35 : std_logic;
    signal l1_single_jet120er2p5 : std_logic;
    signal l1_single_mu0_emtf : std_logic;
    signal l1_single_mu22_bmtf : std_logic;
    signal l1_single_mu22_emtf : std_logic;

-- ========================================================