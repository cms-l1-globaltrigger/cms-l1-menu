-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_0_1

-- Unique ID of L1 Trigger Menu:
-- 88611f82-f9d5-4db8-917c-95d140b6644a

-- Unique ID of firmware implementation:
-- c9eecec0-6ade-4733-b1f9-31711d57aa7c

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.13.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i107 : std_logic;
    signal single_ext_i84 : std_logic;
    signal single_ext_i89 : std_logic;
    signal muon_shower1_i59 : std_logic;
    signal single_htt_i110 : std_logic;
    signal single_eg_i114 : std_logic;
    signal single_jet_i127 : std_logic;
    signal single_mu_i130 : std_logic;
    signal single_mu_i132 : std_logic;
    signal single_mu_i136 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_and_ref4_vme : std_logic;
    signal l1_bptx_not_or_vme : std_logic;
    signal l1_mu_shower_one_tight : std_logic;
    signal l1_first_collision_in_orbit : std_logic;
    signal l1_htt200er : std_logic;
    signal l1_single_eg10er2p5 : std_logic;
    signal l1_single_jet35er2p5 : std_logic;
    signal l1_single_mu0_dq : std_logic;
    signal l1_single_mu0_omtf : std_logic;
    signal l1_single_mu_cosmics_bmtf : std_logic;

-- ========================================================