-- ========================================================
-- from VHDL producer:

-- Module ID: 2

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_1_0

-- Unique ID of L1 Trigger Menu:
-- 11f4244d-31e8-434f-b121-3188fa41b985

-- Unique ID of firmware implementation:
-- c8183b8a-5519-47a4-ad38-1ceb98bede21

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.13.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i86 : std_logic;
    signal single_ext_i91 : std_logic;
    signal muon_shower0_i60 : std_logic;
    signal single_htt_i112 : std_logic;
    signal single_eg_i118 : std_logic;
    signal single_jet_i119 : std_logic;
    signal single_jet_i125 : std_logic;
    signal single_jet_i126 : std_logic;
    signal single_mu_i129 : std_logic;
    signal single_mu_i133 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_beam_gas_b2_vme : std_logic;
    signal l1_bptx_or_ref4_vme : std_logic;
    signal l1_mu_shower_one_nominal : std_logic;
    signal l1_htt360er : std_logic;
    signal l1_single_eg8er2p5 : std_logic;
    signal l1_single_jet120 : std_logic;
    signal l1_single_jet35_fwd3p0 : std_logic;
    signal l1_single_mu0_bmtf : std_logic;
    signal l1_single_mu22 : std_logic;

-- ========================================================