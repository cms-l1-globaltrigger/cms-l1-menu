-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_1_0

-- Unique ID of L1 Trigger Menu:
-- 11f4244d-31e8-434f-b121-3188fa41b985

-- Unique ID of firmware implementation:
-- c8183b8a-5519-47a4-ad38-1ceb98bede21

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.13.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i108 : std_logic;
    signal single_ext_i138 : std_logic;
    signal single_ext_i84 : std_logic;
    signal single_ext_i89 : std_logic;
    signal single_htt_i110 : std_logic;
    signal single_eg_i114 : std_logic;
    signal single_jet_i127 : std_logic;
    signal single_mu_i130 : std_logic;
    signal single_mu_i132 : std_logic;
    signal single_mu_i136 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_and_ref4_vme : std_logic;
    signal l1_bptx_not_or_vme : std_logic;
    signal l1_first_collision_in_train : std_logic;
    signal l1_htt200er : std_logic;
    signal l1_single_eg10er2p5 : std_logic;
    signal l1_single_jet35er2p5 : std_logic;
    signal l1_single_mu0_dq : std_logic;
    signal l1_single_mu0_omtf : std_logic;
    signal l1_single_mu_cosmics_bmtf : std_logic;
    signal l1_unpaired_bunch_bptx_minus : std_logic;

-- ========================================================