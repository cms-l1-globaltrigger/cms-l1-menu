-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2024_v1_0_6

-- Unique ID of L1 Trigger Menu:
-- df279223-6b48-4a59-b67a-2a36dee99794

-- Unique ID of firmware implementation:
-- b76120f9-d3d6-4ba7-bf26-6c1c26c13e0d

-- Scale set:
-- scales_2023_02_16

-- VHDL producer
-- version: 2.20.1
-- hash value: 37aeed0f04da76b667e2567c8eee7fb6e0bbfdcc7e4a47a65d22d7168cf55357

-- tmEventSetup
-- version: 0.13.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i10 : std_logic;
    signal single_ext_i175 : std_logic;
    signal single_ext_i5 : std_logic;
    signal single_etmhf_i35 : std_logic;
    signal single_htt_i177 : std_logic;
    signal single_htt_i180 : std_logic;
    signal double_eg_i166 : std_logic;
    signal double_jet_i170 : std_logic;
    signal single_eg_i186 : std_logic;
    signal single_eg_i245 : std_logic;
    signal single_eg_i249 : std_logic;
    signal single_eg_i253 : std_logic;
    signal single_eg_i46 : std_logic;
    signal single_jet_i49 : std_logic;
    signal single_jet_i50 : std_logic;
    signal single_jet_i51 : std_logic;
    signal single_jet_i54 : std_logic;
    signal single_mu_i59 : std_logic;
    signal single_mu_i60 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_beam_gas_b2_vme : std_logic;
    signal l1_bptx_or_ref4_vme : std_logic;
    signal l1_etmhf100 : std_logic;
    signal l1_htt255er : std_logic;
    signal l1_htt450er : std_logic;
    signal l1_hcal_laser_mon_veto : std_logic;
    signal l1_single_eg26er2p5 : std_logic;
    signal l1_single_eg42er2p5 : std_logic;
    signal l1_double_eg_22_10_er2p5 : std_logic;
    signal l1_single_iso_eg32er2p5 : std_logic;
    signal l1_single_iso_eg34er2p5 : std_logic;
    signal l1_single_jet35er2p5 : std_logic;
    signal l1_single_jet35_fwd3p0 : std_logic;
    signal l1_single_jet120 : std_logic;
    signal l1_double_jet100er2p5 : std_logic;
    signal l1_single_mu0_dq : std_logic;
    signal l1_single_mu0_bmtf : std_logic;
    signal l1_single_iso_eg24er2p1 : std_logic;
    signal l1_single_iso_eg28er2p5 : std_logic;

-- ========================================================