-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2023_v1_1_3

-- Unique ID of L1 Trigger Menu:
-- 4998ea81-aafe-4973-ba76-351aa728a934

-- Unique ID of firmware implementation:
-- 2a223afd-4dc1-482f-9a53-b528d8dc0ac6

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.14.2

-- tmEventSetup version
-- v0.11.2

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i10 : std_logic;
    signal single_ext_i179 : std_logic;
    signal single_ext_i5 : std_logic;
    signal single_ett_i36 : std_logic;
    signal single_htt_i181 : std_logic;
    signal single_htt_i184 : std_logic;
    signal double_eg_i170 : std_logic;
    signal double_jet_i174 : std_logic;
    signal single_eg_i187 : std_logic;
    signal single_eg_i193 : std_logic;
    signal single_eg_i197 : std_logic;
    signal single_eg_i201 : std_logic;
    signal single_eg_i43 : std_logic;
    signal single_eg_i44 : std_logic;
    signal single_jet_i208 : std_logic;
    signal single_jet_i49 : std_logic;
    signal single_jet_i50 : std_logic;
    signal single_mu_i211 : std_logic;
    signal single_mu_i220 : std_logic;
    signal single_mu_i64 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_beam_gas_b2_vme : std_logic;
    signal l1_bptx_or_ref4_vme : std_logic;
    signal l1_ett2000 : std_logic;
    signal l1_single_eg8er2p5 : std_logic;
    signal l1_single_eg10er2p5 : std_logic;
    signal l1_single_jet35_fwd3p0 : std_logic;
    signal l1_single_mu22_bmtf : std_logic;
    signal l1_single_mu_cosmics_omtf : std_logic;
    signal l1_double_eg_22_10_er2p5 : std_logic;
    signal l1_double_jet100er2p5 : std_logic;
    signal l1_hcal_laser_mon_veto : std_logic;
    signal l1_htt255er : std_logic;
    signal l1_htt450er : std_logic;
    signal l1_single_eg36er2p5 : std_logic;
    signal l1_single_iso_eg24er2p1 : std_logic;
    signal l1_single_iso_eg28er2p5 : std_logic;
    signal l1_single_iso_eg32er2p5 : std_logic;
    signal l1_single_jet180 : std_logic;
    signal l1_single_mu18 : std_logic;

-- ========================================================